module abc ();
endmodule
